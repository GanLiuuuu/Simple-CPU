module ALU()
