`timescale 1ns / 1ps

module instruction_fetch(
   input wire clk,             // 时钟信号
   input wire rst,             // 复位信号
   input wire [31:0] PC,       // 程序计数器
   output [31:0] instruction, // 输出指令
   
   //UART
   input upg_rst_i,  // UPG reset (Active High)
   input upg_clk_i,  // UPG clock (10MHz)
   input upg_wen_i,  // UPG write enable
   input [13:0] upg_adr_i,  // UPG write address
   input [31:0] upg_dat_i,  // UPG write data
   input upg_done_i  // 1 if program finished
    );
    
    wire kickOff = upg_rst_i | (~upg_rst_i & upg_done_i);
    prgrom instmesm (
        .clka(kickOff ? clk : upg_clk_i),
        .wea(kickOff ? 1'b0 : upg_wen_i),
        .addra(kickOff ? PC[15:2] : upg_adr_i),
        .dina(kickOff ? 32'h00000000 : upg_dat_i),
        .douta(instruction)
    );

endmodule
